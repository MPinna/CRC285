library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity XOR_LUT is
    generic( Nbit : positive := 8);
    port (
        d_in    : in    std_logic_vector(Nbit - 1 downto 0);
        d_out   : out   std_logic_vector(Nbit - 1 downto 0)
    );
end entity XOR_LUT;

architecture rtl of XOR_LUT is
    
    constant GENERATOR_LEN  :   natural := 8;

    signal  addr_int     :   integer range 0 to 255;
    
    type lut_t is array (0 to 255) of std_logic_vector(GENERATOR_LEN -1 downto 0);
    
    constant lut: lut_t :=
    (
        "00000000", "00011101", "00111010", "00100111", "01110100", "01101001", "01001110", "01010011",
        "11101000", "11110101", "11010010", "11001111", "10011100", "10000001", "10100110", "10111011",
        "11001101", "11010000", "11110111", "11101010", "10111001", "10100100", "10000011", "10011110",
        "00100101", "00111000", "00011111", "00000010", "01010001", "01001100", "01101011", "01110110",
        "10000111", "10011010", "10111101", "10100000", "11110011", "11101110", "11001001", "11010100",
        "01101111", "01110010", "01010101", "01001000", "00011011", "00000110", "00100001", "00111100",
        "01001010", "01010111", "01110000", "01101101", "00111110", "00100011", "00000100", "00011001",
        "10100010", "10111111", "10011000", "10000101", "11010110", "11001011", "11101100", "11110001",
        "00010011", "00001110", "00101001", "00110100", "01100111", "01111010", "01011101", "01000000",
        "11111011", "11100110", "11000001", "11011100", "10001111", "10010010", "10110101", "10101000",
        "11011110", "11000011", "11100100", "11111001", "10101010", "10110111", "10010000", "10001101",
        "00110110", "00101011", "00001100", "00010001", "01000010", "01011111", "01111000", "01100101",
        "10010100", "10001001", "10101110", "10110011", "11100000", "11111101", "11011010", "11000111",
        "01111100", "01100001", "01000110", "01011011", "00001000", "00010101", "00110010", "00101111",
        "01011001", "01000100", "01100011", "01111110", "00101101", "00110000", "00010111", "00001010",
        "10110001", "10101100", "10001011", "10010110", "11000101", "11011000", "11111111", "11100010",
        "00100110", "00111011", "00011100", "00000001", "01010010", "01001111", "01101000", "01110101",
        "11001110", "11010011", "11110100", "11101001", "10111010", "10100111", "10000000", "10011101",
        "11101011", "11110110", "11010001", "11001100", "10011111", "10000010", "10100101", "10111000",
        "00000011", "00011110", "00111001", "00100100", "01110111", "01101010", "01001101", "01010000",
        "10100001", "10111100", "10011011", "10000110", "11010101", "11001000", "11101111", "11110010",
        "01001001", "01010100", "01110011", "01101110", "00111101", "00100000", "00000111", "00011010",
        "01101100", "01110001", "01010110", "01001011", "00011000", "00000101", "00100010", "00111111",
        "10000100", "10011001", "10111110", "10100011", "11110000", "11101101", "11001010", "11010111",
        "00110101", "00101000", "00001111", "00010010", "01000001", "01011100", "01111011", "01100110",
        "11011101", "11000000", "11100111", "11111010", "10101001", "10110100", "10010011", "10001110",
        "11111000", "11100101", "11000010", "11011111", "10001100", "10010001", "10110110", "10101011",
        "00010000", "00001101", "00101010", "00110111", "01100100", "01111001", "01011110", "01000011",
        "10110010", "10101111", "10001000", "10010101", "11000110", "11011011", "11111100", "11100001",
        "01011010", "01000111", "01100000", "01111101", "00101110", "00110011", "00010100", "00001001",
        "01111111", "01100010", "01000101", "01011000", "00001011", "00010110", "00110001", "00101100",
        "10010111", "10001010", "10101101", "10110000", "11100011", "11111110", "11011001", "11000100"
    );
begin
    addr_int    <= TO_INTEGER(unsigned(d_in));
    d_out       <= lut(addr_int);
end architecture rtl;